interface fir_filter_if ();

    bit clk_i;
    bit arstn_i;

endinterface 
